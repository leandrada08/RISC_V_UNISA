module MULT (
    input [31:0] a,
    input [31:0] b,
    output [31:0] product
);
    assign product = a * b;
endmodule
